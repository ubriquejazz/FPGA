---------------------------------------------------------------------------
-- Scattered Pilot Detection
--
-- Scattered Pilot -> k-th sub-carrier in an l-th symbol signal
--
-- k = Kmin + 3 * ( l mod 4 - 1 ) + 12 p 	|| p = 0,1, .. N p - 1 
--											|| k = [Kmin, Kmax]
--											|| l = [0, 67]
-- Kmin = 688; Kmax = 7504 (8K Mode)
-- Kmin = 172; Kmax = 1876 (2K Mode)
--
-- offset 			= Kmin + 3 * ( l mod 4 - 1 ) 			|| l = 0 : 67
-- addr_out(i) 		= offset + addr_int(i) 					|| i = 0 : 568
-- comparacion(i) 	= 1 when addr_out(i) = carrier_indx 	|| i = 0 : 568
--
---------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library WORK;
use WORK.mypackage.all;

entity scatt_detector is
	port (
		clk				: IN 	std_logic;
		reset_n 		: IN  std_logic;
		ce				: IN  std_logic;
		carrier_indx	: IN  std_logic_vector(12 downto 0);	-- k 
		frame_indx		: IN  std_logic_vector(6  downto 0);	-- l
		dispersa		: OUT std_logic
	);
end scatt_detector;


architecture Behavioral of scatt_detector is

	constant Kmin2k 	: std_logic_vector(12 downto 0) := conv_std_logic_vector(172, 13);
	constant Kmin8k 	: std_logic_vector(12 downto 0) := conv_std_logic_vector(688, 13);

	type IndicePilotoDispersa is array(0 to 568) of std_logic_vector(12 downto 0);
	signal addr_out		: IndicePilotoDispersa;	
	signal addr_in		: IndicePilotoDispersa := (
								B"0000000000000" , B"0000000001100" , B"0000000011000" , B"0000000100100" ,
								B"0000000110000" , B"0000000111100" , B"0000001001000" , B"0000001010100" ,
								B"0000001100000" , B"0000001101100" , B"0000001111000" , B"0000010000100" ,
								B"0000010010000" , B"0000010011100" , B"0000010101000" , B"0000010110100" ,
								B"0000011000000" , B"0000011001100" , B"0000011011000" , B"0000011100100" ,
								B"0000011110000" , B"0000011111100" , B"0000100001000" , B"0000100010100" ,
								B"0000100100000" , B"0000100101100" , B"0000100111000" , B"0000101000100" ,
								B"0000101010000" , B"0000101011100" , B"0000101101000" , B"0000101110100" ,
								B"0000110000000" , B"0000110001100" , B"0000110011000" , B"0000110100100" ,
								B"0000110110000" , B"0000110111100" , B"0000111001000" , B"0000111010100" ,
								B"0000111100000" , B"0000111101100" , B"0000111111000" , B"0001000000100" ,
								B"0001000010000" , B"0001000011100" , B"0001000101000" , B"0001000110100" ,
								B"0001001000000" , B"0001001001100" , B"0001001011000" , B"0001001100100" ,
								B"0001001110000" , B"0001001111100" , B"0001010001000" , B"0001010010100" ,
								B"0001010100000" , B"0001010101100" , B"0001010111000" , B"0001011000100" ,
								B"0001011010000" , B"0001011011100" , B"0001011101000" , B"0001011110100" ,
								B"0001100000000" , B"0001100001100" , B"0001100011000" , B"0001100100100" ,
								B"0001100110000" , B"0001100111100" , B"0001101001000" , B"0001101010100" ,
								B"0001101100000" , B"0001101101100" , B"0001101111000" , B"0001110000100" ,
								B"0001110010000" , B"0001110011100" , B"0001110101000" , B"0001110110100" ,
								B"0001111000000" , B"0001111001100" , B"0001111011000" , B"0001111100100" ,
								B"0001111110000" , B"0001111111100" , B"0010000001000" , B"0010000010100" ,
								B"0010000100000" , B"0010000101100" , B"0010000111000" , B"0010001000100" ,
								B"0010001010000" , B"0010001011100" , B"0010001101000" , B"0010001110100" ,
								B"0010010000000" , B"0010010001100" , B"0010010011000" , B"0010010100100" ,
								B"0010010110000" , B"0010010111100" , B"0010011001000" , B"0010011010100" ,
								B"0010011100000" , B"0010011101100" , B"0010011111000" , B"0010100000100" ,
								B"0010100010000" , B"0010100011100" , B"0010100101000" , B"0010100110100" ,
								B"0010101000000" , B"0010101001100" , B"0010101011000" , B"0010101100100" ,
								B"0010101110000" , B"0010101111100" , B"0010110001000" , B"0010110010100" ,
								B"0010110100000" , B"0010110101100" , B"0010110111000" , B"0010111000100" ,
								B"0010111010000" , B"0010111011100" , B"0010111101000" , B"0010111110100" ,
								B"0011000000000" , B"0011000001100" , B"0011000011000" , B"0011000100100" ,
								B"0011000110000" , B"0011000111100" , B"0011001001000" , B"0011001010100" ,
								B"0011001100000" , B"0011001101100" , B"0011001111000" , B"0011010000100" ,
								B"0011010010000" , B"0011010011100" , B"0011010101000" , B"0011010110100" ,
								B"0011011000000" , B"0011011001100" , B"0011011011000" , B"0011011100100" ,
								B"0011011110000" , B"0011011111100" , B"0011100001000" , B"0011100010100" ,
								B"0011100100000" , B"0011100101100" , B"0011100111000" , B"0011101000100" ,
								B"0011101010000" , B"0011101011100" , B"0011101101000" , B"0011101110100" ,
								B"0011110000000" , B"0011110001100" , B"0011110011000" , B"0011110100100" ,
								B"0011110110000" , B"0011110111100" , B"0011111001000" , B"0011111010100" ,
								B"0011111100000" , B"0011111101100" , B"0011111111000" , B"0100000000100" ,
								B"0100000010000" , B"0100000011100" , B"0100000101000" , B"0100000110100" ,
								B"0100001000000" , B"0100001001100" , B"0100001011000" , B"0100001100100" ,
								B"0100001110000" , B"0100001111100" , B"0100010001000" , B"0100010010100" ,
								B"0100010100000" , B"0100010101100" , B"0100010111000" , B"0100011000100" ,
								B"0100011010000" , B"0100011011100" , B"0100011101000" , B"0100011110100" ,
								B"0100100000000" , B"0100100001100" , B"0100100011000" , B"0100100100100" ,
								B"0100100110000" , B"0100100111100" , B"0100101001000" , B"0100101010100" ,
								B"0100101100000" , B"0100101101100" , B"0100101111000" , B"0100110000100" ,
								B"0100110010000" , B"0100110011100" , B"0100110101000" , B"0100110110100" ,
								B"0100111000000" , B"0100111001100" , B"0100111011000" , B"0100111100100" ,
								B"0100111110000" , B"0100111111100" , B"0101000001000" , B"0101000010100" ,
								B"0101000100000" , B"0101000101100" , B"0101000111000" , B"0101001000100" ,
								B"0101001010000" , B"0101001011100" , B"0101001101000" , B"0101001110100" ,
								B"0101010000000" , B"0101010001100" , B"0101010011000" , B"0101010100100" ,
								B"0101010110000" , B"0101010111100" , B"0101011001000" , B"0101011010100" ,
								B"0101011100000" , B"0101011101100" , B"0101011111000" , B"0101100000100" ,
								B"0101100010000" , B"0101100011100" , B"0101100101000" , B"0101100110100" ,
								B"0101101000000" , B"0101101001100" , B"0101101011000" , B"0101101100100" ,
								B"0101101110000" , B"0101101111100" , B"0101110001000" , B"0101110010100" ,
								B"0101110100000" , B"0101110101100" , B"0101110111000" , B"0101111000100" ,
								B"0101111010000" , B"0101111011100" , B"0101111101000" , B"0101111110100" ,
								B"0110000000000" , B"0110000001100" , B"0110000011000" , B"0110000100100" ,
								B"0110000110000" , B"0110000111100" , B"0110001001000" , B"0110001010100" ,
								B"0110001100000" , B"0110001101100" , B"0110001111000" , B"0110010000100" ,
								B"0110010010000" , B"0110010011100" , B"0110010101000" , B"0110010110100" ,
								B"0110011000000" , B"0110011001100" , B"0110011011000" , B"0110011100100" ,
								B"0110011110000" , B"0110011111100" , B"0110100001000" , B"0110100010100" ,
								B"0110100100000" , B"0110100101100" , B"0110100111000" , B"0110101000100" ,
								B"0110101010000" , B"0110101011100" , B"0110101101000" , B"0110101110100" ,
								B"0110110000000" , B"0110110001100" , B"0110110011000" , B"0110110100100" ,
								B"0110110110000" , B"0110110111100" , B"0110111001000" , B"0110111010100" ,
								B"0110111100000" , B"0110111101100" , B"0110111111000" , B"0111000000100" ,
								B"0111000010000" , B"0111000011100" , B"0111000101000" , B"0111000110100" ,
								B"0111001000000" , B"0111001001100" , B"0111001011000" , B"0111001100100" ,
								B"0111001110000" , B"0111001111100" , B"0111010001000" , B"0111010010100" ,
								B"0111010100000" , B"0111010101100" , B"0111010111000" , B"0111011000100" ,
								B"0111011010000" , B"0111011011100" , B"0111011101000" , B"0111011110100" ,
								B"0111100000000" , B"0111100001100" , B"0111100011000" , B"0111100100100" ,
								B"0111100110000" , B"0111100111100" , B"0111101001000" , B"0111101010100" ,
								B"0111101100000" , B"0111101101100" , B"0111101111000" , B"0111110000100" ,
								B"0111110010000" , B"0111110011100" , B"0111110101000" , B"0111110110100" ,
								B"0111111000000" , B"0111111001100" , B"0111111011000" , B"0111111100100" ,
								B"0111111110000" , B"0111111111100" , B"1000000001000" , B"1000000010100" ,
								B"1000000100000" , B"1000000101100" , B"1000000111000" , B"1000001000100" ,
								B"1000001010000" , B"1000001011100" , B"1000001101000" , B"1000001110100" ,
								B"1000010000000" , B"1000010001100" , B"1000010011000" , B"1000010100100" ,
								B"1000010110000" , B"1000010111100" , B"1000011001000" , B"1000011010100" ,
								B"1000011100000" , B"1000011101100" , B"1000011111000" , B"1000100000100" ,
								B"1000100010000" , B"1000100011100" , B"1000100101000" , B"1000100110100" ,
								B"1000101000000" , B"1000101001100" , B"1000101011000" , B"1000101100100" ,
								B"1000101110000" , B"1000101111100" , B"1000110001000" , B"1000110010100" ,
								B"1000110100000" , B"1000110101100" , B"1000110111000" , B"1000111000100" ,
								B"1000111010000" , B"1000111011100" , B"1000111101000" , B"1000111110100" ,
								B"1001000000000" , B"1001000001100" , B"1001000011000" , B"1001000100100" ,
								B"1001000110000" , B"1001000111100" , B"1001001001000" , B"1001001010100" ,
								B"1001001100000" , B"1001001101100" , B"1001001111000" , B"1001010000100" ,
								B"1001010010000" , B"1001010011100" , B"1001010101000" , B"1001010110100" ,
								B"1001011000000" , B"1001011001100" , B"1001011011000" , B"1001011100100" ,
								B"1001011110000" , B"1001011111100" , B"1001100001000" , B"1001100010100" ,
								B"1001100100000" , B"1001100101100" , B"1001100111000" , B"1001101000100" ,
								B"1001101010000" , B"1001101011100" , B"1001101101000" , B"1001101110100" ,
								B"1001110000000" , B"1001110001100" , B"1001110011000" , B"1001110100100" ,
								B"1001110110000" , B"1001110111100" , B"1001111001000" , B"1001111010100" ,
								B"1001111100000" , B"1001111101100" , B"1001111111000" , B"1010000000100" ,
								B"1010000010000" , B"1010000011100" , B"1010000101000" , B"1010000110100" ,
								B"1010001000000" , B"1010001001100" , B"1010001011000" , B"1010001100100" ,
								B"1010001110000" , B"1010001111100" , B"1010010001000" , B"1010010010100" ,
								B"1010010100000" , B"1010010101100" , B"1010010111000" , B"1010011000100" ,
								B"1010011010000" , B"1010011011100" , B"1010011101000" , B"1010011110100" ,
								B"1010100000000" , B"1010100001100" , B"1010100011000" , B"1010100100100" ,
								B"1010100110000" , B"1010100111100" , B"1010101001000" , B"1010101010100" ,
								B"1010101100000" , B"1010101101100" , B"1010101111000" , B"1010110000100" ,
								B"1010110010000" , B"1010110011100" , B"1010110101000" , B"1010110110100" ,
								B"1010111000000" , B"1010111001100" , B"1010111011000" , B"1010111100100" ,
								B"1010111110000" , B"1010111111100" , B"1011000001000" , B"1011000010100" ,
								B"1011000100000" , B"1011000101100" , B"1011000111000" , B"1011001000100" ,
								B"1011001010000" , B"1011001011100" , B"1011001101000" , B"1011001110100" ,
								B"1011010000000" , B"1011010001100" , B"1011010011000" , B"1011010100100" ,
								B"1011010110000" , B"1011010111100" , B"1011011001000" , B"1011011010100" ,
								B"1011011100000" , B"1011011101100" , B"1011011111000" , B"1011100000100" ,
								B"1011100010000" , B"1011100011100" , B"1011100101000" , B"1011100110100" ,
								B"1011101000000" , B"1011101001100" , B"1011101011000" , B"1011101100100" ,
								B"1011101110000" , B"1011101111100" , B"1011110001000" , B"1011110010100" ,
								B"1011110100000" , B"1011110101100" , B"1011110111000" , B"1011111000100" , 
								B"1011111010000" , B"1011111011100" , B"1011111101000" , B"1011111110100" , 
								B"1100000000000" , B"1100000001100" , B"1100000011000" , B"1100000100100" , 
								B"1100000110000" , B"1100000111100" , B"1100001001000" , B"1100001010100" , 
								B"1100001100000" , B"1100001101100" , B"1100001111000" , B"1100010000100" , 
								B"1100010010000" , B"1100010011100" , B"1100010101000" , B"1100010110100" , 
								B"1100011000000" , B"1100011001100" , B"1100011011000" , B"1100011100100" , 
								B"1100011110000" , B"1100011111100" , B"1100100001000" , B"1100100010100" , 
								B"1100100100000" , B"1100100101100" , B"1100100111000" , B"1100101000100" , 
								B"1100101010000" , B"1100101011100" , B"1100101101000" , B"1100101110100" , 
								B"1100110000000" , B"1100110001100" , B"1100110011000" , B"1100110100100" , 
								B"1100110110000" , B"1100110111100" , B"1100111001000" , B"1100111010100" , 
								B"1100111100000" , B"1100111101100" , B"1100111111000" , B"1101000000100" , 
								B"1101000010000" , B"1101000011100" , B"1101000101000" , B"1101000110100" , 
								B"1101001000000" , B"1101001001100" , B"1101001011000" , B"1101001100100" , 
								B"1101001110000" , B"1101001111100" , B"1101010001000" , B"1101010010100" ,
								B"1101010100000" );
											
	COMPONENT scatt_adder
	PORT(
		clk 		: IN 	std_logic;
		reset_n 	: IN 	std_logic;
		ce 			: IN 	std_logic;
		A 			: IN 	std_logic_vector(12 downto 0);
		B 			: IN 	std_logic_vector(12 downto 0);          
		C 			: OUT 	std_logic_vector(12 downto 0)
		);
	END COMPONENT;
	
	COMPONENT scatt_comp
	PORT(
		clk 		: IN 	std_logic;
		reset_n 	: IN 	std_logic;
		ce 			: IN 	std_logic;
		A 			: IN 	std_logic_vector(12 downto 0);
		B 			: IN 	std_logic_vector(12 downto 0);          
		C 			: OUT 	std_logic
		);
	END COMPONENT;

	signal offset2k		: std_logic_vector(12 downto 0);
	signal offset8k		: std_logic_vector(12 downto 0);
	signal comparacion 	: std_logic_vector(568 downto 0);
	
begin

	-- 1� Offset 			ready at	 start0 + 5
	process(clk)
	begin
		if clk'event and clk = '1' then
			if reset_n = '0' then
				offset2k <= (others => '0');
				offset8k <= (others => '0');
			elsif ce = '1' then
				offset2k <= Kmin2k + "11" * frame_indx(1 downto 0);
				offset8k <= Kmin8k + "11" * frame_indx(1 downto 0);
			end if;
		end if;
	end process;

	-- 2� Adders 			ready at	 start0 + 6
	gen_sumadores: for i in 0 to 568 generate
		Inst_sumador: scatt_adder PORT MAP(
			clk 		=> clk,
			reset_n 	=> reset_n,
			ce			=> ce,
			A			=> offset8k,
			B  		=> addr_in(i),
			C 			=> addr_out(i)
		);
	end generate;
		
	-- 3� Comparison	 	ready at	start0 + 7
	gen_comparaciones: for i in 0 to 568 generate
		Inst_comparador: scatt_comp PORT MAP(
			clk 		=> clk,
			reset_n 	=> reset_n,
			ce			=> ce,
			A 			=> addr_out(i),
			B 			=> carrier_indx,	
			C 			=> comparacion(i)
		);
	end generate;
	
	-- 4� Comparison 		ready at	start0 + 8
	process(clk)
	begin
		if clk'event and clk = '1' then
			if reset_n = '0' then
				dispersa <= '0';
			elsif ce = '1' then
				if (comparacion = conv_std_logic_vector(0, 568)) then
					dispersa	<= '0';
				else
					dispersa <= '1';
				end if;	
			end if;
		end if;
	end process;

	--	dispersa  <= '0' when comparacion = conv_std_logic_vector(0, 504) else '1'; 
	
end Behavioral;